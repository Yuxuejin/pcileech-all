//
// PCILeech FPGA.
//
// PCIe BAR PIO controller.
//
// The PCILeech BAR PIO controller allows for easy user-implementation on top
// of the PCILeech AXIS128 PCIe TLP streaming interface.
// The controller consists of a read engine and a write engine and pluggable
// user-implemented PCIe BAR implementations (found at bottom of the file).
//
// Considerations:
// - The core handles 1 DWORD read + 1 DWORD write per CLK max. If a lot of
//   data is written / read from the TLP streaming interface the core may
//   drop packet silently.
// - The core reads 1 DWORD of data (without byte enable) per CLK.
// - The core writes 1 DWORD of data (with byte enable) per CLK.
// - All user-implemented cores must have the same latency in CLKs for the
//   returned read data or else undefined behavior will take place.
// - 32-bit addresses are passed for read/writes. Larger BARs than 4GB are
//   not supported due to addressing constraints. Lower bits (LSBs) are the
//   BAR offset, Higher bits (MSBs) are the 32-bit base address of the BAR.
// - DO NOT edit read/write engines.
// - DO edit pcileech_tlps128_bar_controller (to swap bar implementations).
// - DO edit the bar implementations (at bottom of the file, if neccessary).
//
// Example implementations exists below, swap out any of the example cores
// against a core of your use case, or modify existing cores.
// Following test cores exist (see below in this file):
// - pcileech_bar_impl_zerowrite4k = zero-initialized read/write BAR.
//     It's possible to modify contents by use of .coe file.
// - pcileech_bar_impl_loopaddr = test core that loops back the 32-bit
//     address of the current read. Does not support writes.
// - pcileech_bar_impl_none = core without any reply.
// 
// (c) Ulf Frisk, 2024
// Author: Ulf Frisk, pcileech@frizk.net
//

`timescale 1ns / 1ps
`include "pcileech_header.svh"

module pcileech_tlps128_bar_controller(
    input                   rst,
    input                   clk,
    input                   bar_en,
    input [15:0]            pcie_id,
    input [31:0]            base_address_register,
    IfAXIS128.sink_lite     tlps_in,
    IfAXIS128.source        tlps_out
);
    
    // ------------------------------------------------------------------------
    // 1: TLP RECEIVE:
    // Receive incoming BAR requests from the TLP stream:
    // send them onwards to read and write FIFOs
    // ------------------------------------------------------------------------
    wire in_is_wr_ready;
    bit  in_is_wr_last;
    wire in_is_first    = tlps_in.tuser[0];
    wire in_is_bar      = bar_en && (tlps_in.tuser[8:2] != 0);
    wire in_is_rd       = (in_is_first && tlps_in.tlast && ((tlps_in.tdata[31:25] == 7'b0000000) || (tlps_in.tdata[31:25] == 7'b0010000) || (tlps_in.tdata[31:24] == 8'b00000010)));
    wire in_is_wr       = in_is_wr_last || (in_is_first && in_is_wr_ready && ((tlps_in.tdata[31:25] == 7'b0100000) || (tlps_in.tdata[31:25] == 7'b0110000) || (tlps_in.tdata[31:24] == 8'b01000010)));
    
    always @ ( posedge clk )
        if ( rst ) begin
            in_is_wr_last <= 0;
        end
        else if ( tlps_in.tvalid ) begin
            in_is_wr_last <= !tlps_in.tlast && in_is_wr;
        end
    
    wire [6:0]  wr_bar;
    wire [31:0] wr_addr;
    wire [3:0]  wr_be;
    wire [31:0] wr_data;
    wire        wr_valid;
    wire [87:0] rd_req_ctx;
    wire [6:0]  rd_req_bar;
    wire [31:0] rd_req_addr;
    wire        rd_req_valid;
    wire [87:0] rd_rsp_ctx;
    wire [31:0] rd_rsp_data;
    wire        rd_rsp_valid;
        
    pcileech_tlps128_bar_rdengine i_pcileech_tlps128_bar_rdengine(
        .rst            ( rst                           ),
        .clk            ( clk                           ),
        // TLPs:
        .pcie_id        ( pcie_id                       ),
        .tlps_in        ( tlps_in                       ),
        .tlps_in_valid  ( tlps_in.tvalid && in_is_bar && in_is_rd ),
        .tlps_out       ( tlps_out                      ),
        // BAR reads:
        .rd_req_ctx     ( rd_req_ctx                    ),
        .rd_req_bar     ( rd_req_bar                    ),
        .rd_req_addr    ( rd_req_addr                   ),
        .rd_req_valid   ( rd_req_valid                  ),
        .rd_rsp_ctx     ( rd_rsp_ctx                    ),
        .rd_rsp_data    ( rd_rsp_data                   ),
        .rd_rsp_valid   ( rd_rsp_valid                  )
    );

    pcileech_tlps128_bar_wrengine i_pcileech_tlps128_bar_wrengine(
        .rst            ( rst                           ),
        .clk            ( clk                           ),
        // TLPs:
        .tlps_in        ( tlps_in                       ),
        .tlps_in_valid  ( tlps_in.tvalid && in_is_bar && in_is_wr ),
        .tlps_in_ready  ( in_is_wr_ready                ),
        // outgoing BAR writes:
        .wr_bar         ( wr_bar                        ),
        .wr_addr        ( wr_addr                       ),
        .wr_be          ( wr_be                         ),
        .wr_data        ( wr_data                       ),
        .wr_valid       ( wr_valid                      )
    );
    
    wire [87:0] bar_rsp_ctx[7];
    wire [31:0] bar_rsp_data[7];
    wire        bar_rsp_valid[7];
    
    assign rd_rsp_ctx = bar_rsp_valid[0] ? bar_rsp_ctx[0] :
                        bar_rsp_valid[1] ? bar_rsp_ctx[1] :
                        bar_rsp_valid[2] ? bar_rsp_ctx[2] :
                        bar_rsp_valid[3] ? bar_rsp_ctx[3] :
                        bar_rsp_valid[4] ? bar_rsp_ctx[4] :
                        bar_rsp_valid[5] ? bar_rsp_ctx[5] :
                        bar_rsp_valid[6] ? bar_rsp_ctx[6] : 0;
    assign rd_rsp_data = bar_rsp_valid[0] ? bar_rsp_data[0] :
                        bar_rsp_valid[1] ? bar_rsp_data[1] :
                        bar_rsp_valid[2] ? bar_rsp_data[2] :
                        bar_rsp_valid[3] ? bar_rsp_data[3] :
                        bar_rsp_valid[4] ? bar_rsp_data[4] :
                        bar_rsp_valid[5] ? bar_rsp_data[5] :
                        bar_rsp_valid[6] ? bar_rsp_data[6] : 0;
    assign rd_rsp_valid = bar_rsp_valid[0] || bar_rsp_valid[1] || bar_rsp_valid[2] || bar_rsp_valid[3] || bar_rsp_valid[4] || bar_rsp_valid[5] || bar_rsp_valid[6];
    
    pcileech_bar_impl_ar9287_wifi i_bar0(
        .rst                   ( rst                           ),
        .clk                   ( clk                           ),
        .wr_addr               ( wr_addr                       ),
        .wr_be                 ( wr_be                         ),
        .wr_data               ( wr_data                       ),
        .wr_valid              ( wr_valid && wr_bar[0]         ),
        .rd_req_ctx            ( rd_req_ctx                    ),
        .rd_req_addr           ( rd_req_addr                   ),
        .rd_req_valid          ( rd_req_valid && rd_req_bar[0] ),
        .base_address_register ( base_address_register         ),
        .rd_rsp_ctx            ( bar_rsp_ctx[0]                ),
        .rd_rsp_data           ( bar_rsp_data[0]               ),
        .rd_rsp_valid          ( bar_rsp_valid[0]              )
    );
    
    pcileech_bar_impl_loopaddr i_bar1(
        .rst            ( rst                           ),
        .clk            ( clk                           ),
        .wr_addr        ( wr_addr                       ),
        .wr_be          ( wr_be                         ),
        .wr_data        ( wr_data                       ),
        .wr_valid       ( wr_valid && wr_bar[1]         ),
        .rd_req_ctx     ( rd_req_ctx                    ),
        .rd_req_addr    ( rd_req_addr                   ),
        .rd_req_valid   ( rd_req_valid && rd_req_bar[1] ),
        .rd_rsp_ctx     ( bar_rsp_ctx[1]                ),
        .rd_rsp_data    ( bar_rsp_data[1]               ),
        .rd_rsp_valid   ( bar_rsp_valid[1]              )
    );
    
    pcileech_bar_impl_none i_bar2(
        .rst            ( rst                           ),
        .clk            ( clk                           ),
        .wr_addr        ( wr_addr                       ),
        .wr_be          ( wr_be                         ),
        .wr_data        ( wr_data                       ),
        .wr_valid       ( wr_valid && wr_bar[2]         ),
        .rd_req_ctx     ( rd_req_ctx                    ),
        .rd_req_addr    ( rd_req_addr                   ),
        .rd_req_valid   ( rd_req_valid && rd_req_bar[2] ),
        .rd_rsp_ctx     ( bar_rsp_ctx[2]                ),
        .rd_rsp_data    ( bar_rsp_data[2]               ),
        .rd_rsp_valid   ( bar_rsp_valid[2]              )
    );
    
    pcileech_bar_impl_none i_bar3(
        .rst            ( rst                           ),
        .clk            ( clk                           ),
        .wr_addr        ( wr_addr                       ),
        .wr_be          ( wr_be                         ),
        .wr_data        ( wr_data                       ),
        .wr_valid       ( wr_valid && wr_bar[3]         ),
        .rd_req_ctx     ( rd_req_ctx                    ),
        .rd_req_addr    ( rd_req_addr                   ),
        .rd_req_valid   ( rd_req_valid && rd_req_bar[3] ),
        .rd_rsp_ctx     ( bar_rsp_ctx[3]                ),
        .rd_rsp_data    ( bar_rsp_data[3]               ),
        .rd_rsp_valid   ( bar_rsp_valid[3]              )
    );
    
    pcileech_bar_impl_none i_bar4(
        .rst            ( rst                           ),
        .clk            ( clk                           ),
        .wr_addr        ( wr_addr                       ),
        .wr_be          ( wr_be                         ),
        .wr_data        ( wr_data                       ),
        .wr_valid       ( wr_valid && wr_bar[4]         ),
        .rd_req_ctx     ( rd_req_ctx                    ),
        .rd_req_addr    ( rd_req_addr                   ),
        .rd_req_valid   ( rd_req_valid && rd_req_bar[4] ),
        .rd_rsp_ctx     ( bar_rsp_ctx[4]                ),
        .rd_rsp_data    ( bar_rsp_data[4]               ),
        .rd_rsp_valid   ( bar_rsp_valid[4]              )
    );
    
    pcileech_bar_impl_none i_bar5(
        .rst            ( rst                           ),
        .clk            ( clk                           ),
        .wr_addr        ( wr_addr                       ),
        .wr_be          ( wr_be                         ),
        .wr_data        ( wr_data                       ),
        .wr_valid       ( wr_valid && wr_bar[5]         ),
        .rd_req_ctx     ( rd_req_ctx                    ),
        .rd_req_addr    ( rd_req_addr                   ),
        .rd_req_valid   ( rd_req_valid && rd_req_bar[5] ),
        .rd_rsp_ctx     ( bar_rsp_ctx[5]                ),
        .rd_rsp_data    ( bar_rsp_data[5]               ),
        .rd_rsp_valid   ( bar_rsp_valid[5]              )
    );
    
    pcileech_bar_impl_none i_bar6_optrom(
        .rst            ( rst                           ),
        .clk            ( clk                           ),
        .wr_addr        ( wr_addr                       ),
        .wr_be          ( wr_be                         ),
        .wr_data        ( wr_data                       ),
        .wr_valid       ( wr_valid && wr_bar[6]         ),
        .rd_req_ctx     ( rd_req_ctx                    ),
        .rd_req_addr    ( rd_req_addr                   ),
        .rd_req_valid   ( rd_req_valid && rd_req_bar[6] ),
        .rd_rsp_ctx     ( bar_rsp_ctx[6]                ),
        .rd_rsp_data    ( bar_rsp_data[6]               ),
        .rd_rsp_valid   ( bar_rsp_valid[6]              )
    );


endmodule



// ------------------------------------------------------------------------
// BAR WRITE ENGINE:
// Receives BAR WRITE TLPs and output BAR WRITE requests.
// Holds a 2048-byte buffer.
// Input flow rate is 16bytes/CLK (max).
// Output flow rate is 4bytes/CLK.
// If write engine overflows incoming TLP is completely discarded silently.
// ------------------------------------------------------------------------
module pcileech_tlps128_bar_wrengine(
    input                   rst,    
    input                   clk,
    // TLPs:
    IfAXIS128.sink_lite     tlps_in,
    input                   tlps_in_valid,
    output                  tlps_in_ready,
    // outgoing BAR writes:
    output bit [6:0]        wr_bar,
    output bit [31:0]       wr_addr,
    output bit [3:0]        wr_be,
    output bit [31:0]       wr_data,
    output bit              wr_valid
);

    wire            f_rd_en;
    wire [127:0]    f_tdata;
    wire [3:0]      f_tkeepdw;
    wire [8:0]      f_tuser;
    wire            f_tvalid;
    
    bit [127:0]     tdata;
    bit [3:0]       tkeepdw;
    bit             tlast;
    
    bit [3:0]       be_first;
    bit [3:0]       be_last;
    bit             first_dw;
    bit [31:0]      addr;

    fifo_141_141_clk1_bar_wr i_fifo_141_141_clk1_bar_wr(
        .srst           ( rst                           ),
        .clk            ( clk                           ),
        .wr_en          ( tlps_in_valid                 ),
        .din            ( {tlps_in.tuser[8:0], tlps_in.tkeepdw, tlps_in.tdata} ),
        .full           (                               ),
        .prog_empty     ( tlps_in_ready                 ),
        .rd_en          ( f_rd_en                       ),
        .dout           ( {f_tuser, f_tkeepdw, f_tdata} ),    
        .empty          (                               ),
        .valid          ( f_tvalid                      )
    );
    
    // STATE MACHINE:
    `define S_ENGINE_IDLE        3'h0
    `define S_ENGINE_FIRST       3'h1
    `define S_ENGINE_4DW_REQDATA 3'h2
    `define S_ENGINE_TX0         3'h4
    `define S_ENGINE_TX1         3'h5
    `define S_ENGINE_TX2         3'h6
    `define S_ENGINE_TX3         3'h7
    (* KEEP = "TRUE" *) bit [3:0] state = `S_ENGINE_IDLE;
    
    assign f_rd_en = (state == `S_ENGINE_IDLE) ||
                     (state == `S_ENGINE_4DW_REQDATA) ||
                     (state == `S_ENGINE_TX3) ||
                     ((state == `S_ENGINE_TX2 && !tkeepdw[3])) ||
                     ((state == `S_ENGINE_TX1 && !tkeepdw[2])) ||
                     ((state == `S_ENGINE_TX0 && !f_tkeepdw[1]));

    always @ ( posedge clk ) begin
        wr_addr     <= addr;
        wr_valid    <= ((state == `S_ENGINE_TX0) && f_tvalid) || (state == `S_ENGINE_TX1) || (state == `S_ENGINE_TX2) || (state == `S_ENGINE_TX3);
        
    end

    always @ ( posedge clk )
        if ( rst ) begin
            state <= `S_ENGINE_IDLE;
        end
        else case ( state )
            `S_ENGINE_IDLE: begin
                state   <= `S_ENGINE_FIRST;
            end
            `S_ENGINE_FIRST: begin
                if ( f_tvalid && f_tuser[0] ) begin
                    wr_bar      <= f_tuser[8:2];
                    tdata       <= f_tdata;
                    tkeepdw     <= f_tkeepdw;
                    tlast       <= f_tuser[1];
                    first_dw    <= 1;
                    be_first    <= f_tdata[35:32];
                    be_last     <= f_tdata[39:36];
                    if ( f_tdata[31:29] == 8'b010 ) begin       // 3 DW header, with data
                        addr    <= { f_tdata[95:66], 2'b00 };
                        state   <= `S_ENGINE_TX3;
                    end
                    else if ( f_tdata[31:29] == 8'b011 ) begin  // 4 DW header, with data
                        addr    <= { f_tdata[127:98], 2'b00 };
                        state   <= `S_ENGINE_4DW_REQDATA;
                    end 
                end
                else begin
                    state   <= `S_ENGINE_IDLE;
                end
            end 
            `S_ENGINE_4DW_REQDATA: begin
                state   <= `S_ENGINE_TX0;
            end
            `S_ENGINE_TX0: begin
                tdata       <= f_tdata;
                tkeepdw     <= f_tkeepdw;
                tlast       <= f_tuser[1];
                addr        <= addr + 4;
                wr_data     <= { f_tdata[0+00+:8], f_tdata[0+08+:8], f_tdata[0+16+:8], f_tdata[0+24+:8] };
                first_dw    <= 0;
                wr_be       <= first_dw ? be_first : (f_tkeepdw[1] ? 4'hf : be_last);
                state       <= f_tvalid ? (f_tkeepdw[1] ? `S_ENGINE_TX1 : `S_ENGINE_FIRST) : `S_ENGINE_IDLE;
            end
            `S_ENGINE_TX1: begin
                addr        <= addr + 4;
                wr_data     <= { tdata[32+00+:8], tdata[32+08+:8], tdata[32+16+:8], tdata[32+24+:8] };
                first_dw    <= 0;
                wr_be       <= first_dw ? be_first : (tkeepdw[2] ? 4'hf : be_last);
                state       <= tkeepdw[2] ? `S_ENGINE_TX2 : `S_ENGINE_FIRST;
            end
            `S_ENGINE_TX2: begin
                addr        <= addr + 4;
                wr_data     <= { tdata[64+00+:8], tdata[64+08+:8], tdata[64+16+:8], tdata[64+24+:8] };
                first_dw    <= 0;
                wr_be       <= first_dw ? be_first : (tkeepdw[3] ? 4'hf : be_last);
                state       <= tkeepdw[3] ? `S_ENGINE_TX3 : `S_ENGINE_FIRST;
            end
            `S_ENGINE_TX3: begin
                addr        <= addr + 4;
                wr_data     <= { tdata[96+00+:8], tdata[96+08+:8], tdata[96+16+:8], tdata[96+24+:8] };
                first_dw    <= 0;
                wr_be       <= first_dw ? be_first : (!tlast ? 4'hf : be_last);
                state       <= !tlast ? `S_ENGINE_TX0 : `S_ENGINE_FIRST;
            end
        endcase

endmodule



// ------------------------------------------------------------------------
// BAR READ ENGINE:
// Receives BAR READ TLPs and output BAR READ requests.
// ------------------------------------------------------------------------
module pcileech_tlps128_bar_rdengine(
    input                   rst,    
    input                   clk,
    // TLPs:
    input [15:0]            pcie_id,
    IfAXIS128.sink_lite     tlps_in,
    input                   tlps_in_valid,
    IfAXIS128.source        tlps_out,
    // BAR reads:
    output [87:0]           rd_req_ctx,
    output [6:0]            rd_req_bar,
    output [31:0]           rd_req_addr,
    output                  rd_req_valid,
    input  [87:0]           rd_rsp_ctx,
    input  [31:0]           rd_rsp_data,
    input                   rd_rsp_valid
);

    // ------------------------------------------------------------------------
    // 1: PROCESS AND QUEUE INCOMING READ TLPs:
    // ------------------------------------------------------------------------
    wire [10:0] rd1_in_dwlen    = (tlps_in.tdata[9:0] == 0) ? 11'd1024 : {1'b0, tlps_in.tdata[9:0]};
    wire [6:0]  rd1_in_bar      = tlps_in.tuser[8:2];
    wire [15:0] rd1_in_reqid    = tlps_in.tdata[63:48];
    wire [7:0]  rd1_in_tag      = tlps_in.tdata[47:40];
    wire [31:0] rd1_in_addr     = { ((tlps_in.tdata[31:29] == 3'b000) ? tlps_in.tdata[95:66] : tlps_in.tdata[127:98]), 2'b00 };
    wire [73:0] rd1_in_data;
    assign rd1_in_data[73:63]   = rd1_in_dwlen;
    assign rd1_in_data[62:56]   = rd1_in_bar;   
    assign rd1_in_data[55:48]   = rd1_in_tag;
    assign rd1_in_data[47:32]   = rd1_in_reqid;
    assign rd1_in_data[31:0]    = rd1_in_addr;
    
    wire        rd1_out_rden;
    wire [73:0] rd1_out_data;
    wire        rd1_out_valid;
    
    fifo_74_74_clk1_bar_rd1 i_fifo_74_74_clk1_bar_rd1(
        .srst           ( rst                           ),
        .clk            ( clk                           ),
        .wr_en          ( tlps_in_valid                 ),
        .din            ( rd1_in_data                   ),
        .full           (                               ),
        .rd_en          ( rd1_out_rden                  ),
        .dout           ( rd1_out_data                  ),    
        .empty          (                               ),
        .valid          ( rd1_out_valid                 )
    );
    
    // ------------------------------------------------------------------------
    // 2: PROCESS AND SPLIT READ TLPs INTO RESPONSE TLP READ REQUESTS AND QUEUE:
    //    (READ REQUESTS LARGER THAN 128-BYTES WILL BE SPLIT INTO MULTIPLE).
    // ------------------------------------------------------------------------
    
    wire [10:0] rd1_out_dwlen       = rd1_out_data[73:63];
    wire [4:0]  rd1_out_dwlen5      = rd1_out_data[67:63];
    wire [4:0]  rd1_out_addr5       = rd1_out_data[6:2];
    
    // 1st "instant" packet:
    wire [4:0]  rd2_pkt1_dwlen_pre  = ((rd1_out_addr5 + rd1_out_dwlen5 > 6'h20) || ((rd1_out_addr5 != 0) && (rd1_out_dwlen5 == 0))) ? (6'h20 - rd1_out_addr5) : rd1_out_dwlen5;
    wire [5:0]  rd2_pkt1_dwlen      = (rd2_pkt1_dwlen_pre == 0) ? 6'h20 : rd2_pkt1_dwlen_pre;
    wire [10:0] rd2_pkt1_dwlen_next = rd1_out_dwlen - rd2_pkt1_dwlen;
    wire        rd2_pkt1_large      = (rd1_out_dwlen > 32) || (rd1_out_dwlen != rd2_pkt1_dwlen);
    wire        rd2_pkt1_tiny       = (rd1_out_dwlen == 1);
    wire [11:0] rd2_pkt1_bc         = rd1_out_dwlen << 2;
    wire [85:0] rd2_pkt1;
    assign      rd2_pkt1[85:74]     = rd2_pkt1_bc;
    assign      rd2_pkt1[73:63]     = rd2_pkt1_dwlen;
    assign      rd2_pkt1[62:0]      = rd1_out_data[62:0];
    
    // Nth packet (if split should take place):
    bit  [10:0] rd2_total_dwlen;
    wire [10:0] rd2_total_dwlen_next = rd2_total_dwlen - 11'h20;
    
    bit  [85:0] rd2_pkt2;
    wire [10:0] rd2_pkt2_dwlen = rd2_pkt2[73:63];
    wire        rd2_pkt2_large = (rd2_total_dwlen > 11'h20);
    
    wire        rd2_out_rden;
    
    // STATE MACHINE:
    `define S2_ENGINE_REQDATA     1'h0
    `define S2_ENGINE_PROCESSING  1'h1
    (* KEEP = "TRUE" *) bit [0:0] state2 = `S2_ENGINE_REQDATA;
    
    always @ ( posedge clk )
        if ( rst ) begin
            state2 <= `S2_ENGINE_REQDATA;
        end
        else case ( state2 )
            `S2_ENGINE_REQDATA: begin
                if ( rd1_out_valid && rd2_pkt1_large ) begin
                    rd2_total_dwlen <= rd2_pkt1_dwlen_next;                             // dwlen (total remaining)
                    rd2_pkt2[85:74] <= rd2_pkt1_dwlen_next << 2;                        // byte-count
                    rd2_pkt2[73:63] <= (rd2_pkt1_dwlen_next > 11'h20) ? 11'h20 : rd2_pkt1_dwlen_next;   // dwlen next
                    rd2_pkt2[62:12] <= rd1_out_data[62:12];                             // various data
                    rd2_pkt2[11:0]  <= rd1_out_data[11:0] + (rd2_pkt1_dwlen << 2);      // base address (within 4k page)
                    state2 <= `S2_ENGINE_PROCESSING;
                end
            end
            `S2_ENGINE_PROCESSING: begin
                if ( rd2_out_rden ) begin
                    rd2_total_dwlen <= rd2_total_dwlen_next;                                // dwlen (total remaining)
                    rd2_pkt2[85:74] <= rd2_total_dwlen_next << 2;                           // byte-count
                    rd2_pkt2[73:63] <= (rd2_total_dwlen_next > 11'h20) ? 11'h20 : rd2_total_dwlen_next;   // dwlen next
                    rd2_pkt2[62:12] <= rd2_pkt2[62:12];                                     // various data
                    rd2_pkt2[11:0]  <= rd2_pkt2[11:0] + (rd2_pkt2_dwlen << 2);              // base address (within 4k page)
                    if ( !rd2_pkt2_large ) begin
                        state2 <= `S2_ENGINE_REQDATA;
                    end
                end
            end
        endcase
    
    assign rd1_out_rden = rd2_out_rden && (((state2 == `S2_ENGINE_REQDATA) && (!rd1_out_valid || rd2_pkt1_tiny)) || ((state2 == `S2_ENGINE_PROCESSING) && !rd2_pkt2_large));

    wire [85:0] rd2_in_data  = (state2 == `S2_ENGINE_REQDATA) ? rd2_pkt1 : rd2_pkt2;
    wire        rd2_in_valid = rd1_out_valid || ((state2 == `S2_ENGINE_PROCESSING) && rd2_out_rden);

    bit  [85:0] rd2_out_data;
    bit         rd2_out_valid;
    always @ ( posedge clk ) begin
        rd2_out_data    <= rd2_in_valid ? rd2_in_data : rd2_out_data;
        rd2_out_valid   <= rd2_in_valid && !rst;
    end

    // ------------------------------------------------------------------------
    // 3: PROCESS EACH READ REQUEST PACKAGE PER INDIVIDUAL 32-bit READ DWORDS:
    // ------------------------------------------------------------------------

    wire [4:0]  rd2_out_dwlen   = rd2_out_data[67:63];
    wire        rd2_out_last    = (rd2_out_dwlen == 1);
    wire [9:0]  rd2_out_dwaddr  = rd2_out_data[11:2];
    
    wire        rd3_enable;
    
    bit         rd3_process_valid;
    bit         rd3_process_first;
    bit         rd3_process_last;
    bit [4:0]   rd3_process_dwlen;
    bit [9:0]   rd3_process_dwaddr;
    bit [85:0]  rd3_process_data;
    wire        rd3_process_next_last = (rd3_process_dwlen == 2);
    wire        rd3_process_nextnext_last = (rd3_process_dwlen <= 3);
    
    assign rd_req_ctx   = { rd3_process_first, rd3_process_last, rd3_process_data };
    assign rd_req_bar   = rd3_process_data[62:56];
    assign rd_req_addr  = { rd3_process_data[31:12], rd3_process_dwaddr, 2'b00 };
    assign rd_req_valid = rd3_process_valid;
    
    // STATE MACHINE:
    `define S3_ENGINE_REQDATA     1'h0
    `define S3_ENGINE_PROCESSING  1'h1
    (* KEEP = "TRUE" *) bit [0:0] state3 = `S3_ENGINE_REQDATA;
    
    always @ ( posedge clk )
        if ( rst ) begin
            rd3_process_valid   <= 1'b0;
            state3              <= `S3_ENGINE_REQDATA;
        end
        else case ( state3 )
            `S3_ENGINE_REQDATA: begin
                if ( rd2_out_valid ) begin
                    rd3_process_valid       <= 1'b1;
                    rd3_process_first       <= 1'b1;                    // FIRST
                    rd3_process_last        <= rd2_out_last;            // LAST (low 5 bits of dwlen == 1, [max pktlen = 0x20))
                    rd3_process_dwlen       <= rd2_out_dwlen;           // PKT LENGTH IN DW
                    rd3_process_dwaddr      <= rd2_out_dwaddr;          // DWADDR OF THIS DWORD
                    rd3_process_data[85:0]  <= rd2_out_data[85:0];      // FORWARD / SAVE DATA
                    if ( !rd2_out_last ) begin
                        state3 <= `S3_ENGINE_PROCESSING;
                    end
                end
                else begin
                    rd3_process_valid       <= 1'b0;
                end
            end
            `S3_ENGINE_PROCESSING: begin
                rd3_process_first           <= 1'b0;                    // FIRST
                rd3_process_last            <= rd3_process_next_last;   // LAST
                rd3_process_dwlen           <= rd3_process_dwlen - 1;   // LEN DEC
                rd3_process_dwaddr          <= rd3_process_dwaddr + 1;  // ADDR INC
                if ( rd3_process_next_last ) begin
                    state3 <= `S3_ENGINE_REQDATA;
                end
            end
        endcase

    assign rd2_out_rden = rd3_enable && (
        ((state3 == `S3_ENGINE_REQDATA) && (!rd2_out_valid || rd2_out_last)) ||
        ((state3 == `S3_ENGINE_PROCESSING) && rd3_process_nextnext_last));
    
    // ------------------------------------------------------------------------
    // 4: PROCESS RESPONSES:
    // ------------------------------------------------------------------------
    
    wire        rd_rsp_first    = rd_rsp_ctx[87];
    wire        rd_rsp_last     = rd_rsp_ctx[86];
    
    wire [9:0]  rd_rsp_dwlen    = rd_rsp_ctx[72:63];
    wire [11:0] rd_rsp_bc       = rd_rsp_ctx[85:74];
    wire [15:0] rd_rsp_reqid    = rd_rsp_ctx[47:32];
    wire [7:0]  rd_rsp_tag      = rd_rsp_ctx[55:48];
    wire [6:0]  rd_rsp_lowaddr  = rd_rsp_ctx[6:0];
    wire [31:0] rd_rsp_addr     = rd_rsp_ctx[31:0];
    wire [31:0] rd_rsp_data_bs  = { rd_rsp_data[7:0], rd_rsp_data[15:8], rd_rsp_data[23:16], rd_rsp_data[31:24] };
    
    // 1: 32-bit -> 128-bit state machine:
    bit [127:0] tdata;
    bit [3:0]   tkeepdw = 0;
    bit         tlast;
    bit         first   = 1;
    wire        tvalid  = tlast || tkeepdw[3];
    
    always @ ( posedge clk )
        if ( rst ) begin
            tkeepdw <= 0;
            tlast   <= 0;
            first   <= 0;
        end
        else if ( rd_rsp_valid && rd_rsp_first ) begin
            tkeepdw         <= 4'b1111;
            tlast           <= rd_rsp_last;
            first           <= 1'b1;
            tdata[31:0]     <= { 22'b0100101000000000000000, rd_rsp_dwlen };            // format, type, length
            tdata[63:32]    <= { pcie_id[7:0], pcie_id[15:8], 4'b0, rd_rsp_bc };        // pcie_id, byte_count
            tdata[95:64]    <= { rd_rsp_reqid, rd_rsp_tag, 1'b0, rd_rsp_lowaddr };      // req_id, tag, lower_addr
            tdata[127:96]   <= rd_rsp_data_bs;
        end
        else begin
            tlast   <= rd_rsp_valid && rd_rsp_last;
            tkeepdw <= tvalid ? (rd_rsp_valid ? 4'b0001 : 4'b0000) : (rd_rsp_valid ? ((tkeepdw << 1) | 1'b1) : tkeepdw);
            first   <= 0;
            if ( rd_rsp_valid ) begin
                if ( tvalid || !tkeepdw[0] )
                    tdata[31:0]   <= rd_rsp_data_bs;
                if ( !tkeepdw[1] )
                    tdata[63:32]  <= rd_rsp_data_bs;
                if ( !tkeepdw[2] )
                    tdata[95:64]  <= rd_rsp_data_bs;
                if ( !tkeepdw[3] )
                    tdata[127:96] <= rd_rsp_data_bs;   
            end
        end
    
    // 2.1 - submit to output fifo - will feed into mux/pcie core.
    fifo_134_134_clk1_bar_rdrsp i_fifo_134_134_clk1_bar_rdrsp(
        .srst           ( rst                       ),
        .clk            ( clk                       ),
        .din            ( { first, tlast, tkeepdw, tdata } ),
        .wr_en          ( tvalid                    ),
        .rd_en          ( tlps_out.tready           ),
        .dout           ( { tlps_out.tuser[0], tlps_out.tlast, tlps_out.tkeepdw, tlps_out.tdata } ),
        .full           (                           ),
        .empty          (                           ),
        .prog_empty     ( rd3_enable                ),
        .valid          ( tlps_out.tvalid           )
    );
    
    assign tlps_out.tuser[1] = tlps_out.tlast;
    assign tlps_out.tuser[8:2] = 0;
    
    // 2.2 - packet count:
    bit [10:0]  pkt_count       = 0;
    wire        pkt_count_dec   = tlps_out.tvalid && tlps_out.tlast;
    wire        pkt_count_inc   = tvalid && tlast;
    wire [10:0] pkt_count_next  = pkt_count + pkt_count_inc - pkt_count_dec;
    assign tlps_out.has_data    = (pkt_count_next > 0);
    
    always @ ( posedge clk ) begin
        pkt_count <= rst ? 0 : pkt_count_next;
    end

endmodule



// ------------------------------------------------------------------------
// Example BAR implementation that does nothing but drop any read/writes
// silently without generating a response.
// This is only recommended for placeholder designs.
// Latency = N/A.
// ------------------------------------------------------------------------
module pcileech_bar_impl_none(
    input               rst,
    input               clk,
    // incoming BAR writes:
    input [31:0]        wr_addr,
    input [3:0]         wr_be,
    input [31:0]        wr_data,
    input               wr_valid,
    // incoming BAR reads:
    input  [87:0]       rd_req_ctx,
    input  [31:0]       rd_req_addr,
    input               rd_req_valid,
    // outgoing BAR read replies:
    output bit [87:0]   rd_rsp_ctx,
    output bit [31:0]   rd_rsp_data,
    output bit          rd_rsp_valid
);

    initial rd_rsp_ctx = 0;
    initial rd_rsp_data = 0;
    initial rd_rsp_valid = 0;

endmodule



// ------------------------------------------------------------------------
// Example BAR implementation of "address loopback" which can be useful
// for testing. Any read to a specific BAR address will result in the
// address as response.
// Latency = 2CLKs.
// ------------------------------------------------------------------------
module pcileech_bar_impl_loopaddr(
    input               rst,
    input               clk,
    // incoming BAR writes:
    input [31:0]        wr_addr,
    input [3:0]         wr_be,
    input [31:0]        wr_data,
    input               wr_valid,
    // incoming BAR reads:
    input [87:0]        rd_req_ctx,
    input [31:0]        rd_req_addr,
    input               rd_req_valid,
    // outgoing BAR read replies:
    output bit [87:0]   rd_rsp_ctx,
    output bit [31:0]   rd_rsp_data,
    output bit          rd_rsp_valid
);

    bit [87:0]      rd_req_ctx_1;
    bit [31:0]      rd_req_addr_1;
    bit             rd_req_valid_1;
    
    always @ ( posedge clk ) begin
        rd_req_ctx_1    <= rd_req_ctx;
        rd_req_addr_1   <= rd_req_addr;
        rd_req_valid_1  <= rd_req_valid;
        rd_rsp_ctx      <= rd_req_ctx_1;
        rd_rsp_data     <= rd_req_addr_1;
        rd_rsp_valid    <= rd_req_valid_1;
    end    

endmodule



// ------------------------------------------------------------------------
// Example BAR implementation of a 4kB writable initial-zero BAR.
// Latency = 2CLKs.
// ------------------------------------------------------------------------
module pcileech_bar_impl_zerowrite4k(
    input               rst,
    input               clk,
    // incoming BAR writes:
    input [31:0]        wr_addr,
    input [3:0]         wr_be,
    input [31:0]        wr_data,
    input               wr_valid,
    // incoming BAR reads:
    input  [87:0]       rd_req_ctx,
    input  [31:0]       rd_req_addr,
    input               rd_req_valid,
    // outgoing BAR read replies:
    output bit [87:0]   rd_rsp_ctx,
    output bit [31:0]   rd_rsp_data,
    output bit          rd_rsp_valid
);

    bit [87:0]  drd_req_ctx;
    bit         drd_req_valid;
    wire [31:0] doutb;
    
    always @ ( posedge clk ) begin
        drd_req_ctx     <= rd_req_ctx;
        drd_req_valid   <= rd_req_valid;
        rd_rsp_ctx      <= drd_req_ctx;
        rd_rsp_valid    <= drd_req_valid;
        rd_rsp_data     <= doutb; 
    end
    
    bram_bar_zero4k i_bram_bar_zero4k(
        // Port A - write:
        .addra  ( wr_addr[11:2]     ),
        .clka   ( clk               ),
        .dina   ( wr_data           ),
        .ena    ( wr_valid          ),
        .wea    ( wr_be             ),
        // Port A - read (2 CLK latency):
        .addrb  ( rd_req_addr[11:2] ),
        .clkb   ( clk               ),
        .doutb  ( doutb             ),
        .enb    ( rd_req_valid      )
    );

endmodule



// ------------------------------------------------------------------------
// pcileech wifi BAR implementation
// Works with Qualcomm Atheros AR9287 chip wifi adapters
// ------------------------------------------------------------------------
module pcileech_bar_impl_ar9287_wifi(
    input               rst,
    input               clk,
    // incoming BAR writes:
    input [31:0]        wr_addr,
    input [3:0]         wr_be,
    input [31:0]        wr_data,
    input               wr_valid,
    // incoming BAR reads:
    input  [87:0]       rd_req_ctx,
    input  [31:0]       rd_req_addr,
    input               rd_req_valid,
    input  [31:0]       base_address_register,
    // outgoing BAR read replies:
    output bit [87:0]   rd_rsp_ctx,
    output bit [31:0]   rd_rsp_data,
    output bit          rd_rsp_valid
);

    bit [87:0]      drd_req_ctx;
    bit [31:0]      drd_req_addr;
    bit             drd_req_valid;

    bit [31:0]      dwr_addr;
    bit [31:0]      dwr_data;
    bit             dwr_valid;

    bit [31:0]      data_32;

    time number = 0;
    
    // 添加统计信息和状态寄存器
    reg [31:0] rx_packets = 0;
    reg [31:0] tx_packets = 0;
    reg [31:0] rx_bytes = 0;
    reg [31:0] tx_bytes = 0;
    reg [31:0] rx_errors = 0;
    reg [31:0] tx_errors = 0;
    reg [3:0] device_state = 0;
    reg [3:0] device_temperature = 4;
    reg [3:0] signal_strength = 0;
    reg [1:0] link_status = 0;
    
    // 添加中断相关寄存器
    reg [31:0] int_status = 0;        // 中断状态寄存器
    reg [31:0] int_mask = 32'hFFFFFFFF; // 中断掩码寄存器，默认全部启用
    reg [31:0] int_cause = 0;         // 中断原因寄存器
    reg [31:0] int_ack = 0;           // 中断确认寄存器
    
    // MSI-X中断表和PBA区域
    reg [127:0] msix_table[16];       // 16个MSI-X表项，每项128位
    reg [31:0] msix_pba = 0;          // Pending Bit Array
    
    // 中断位定义
    localparam INT_RX_COMPLETE = 32'h00000001;  // 接收完成中断
    localparam INT_TX_COMPLETE = 32'h00000002;  // 发送完成中断
    localparam INT_RX_ERROR = 32'h00000004;     // 接收错误中断
    localparam INT_TX_ERROR = 32'h00000008;     // 发送错误中断
    localparam INT_LINK_CHANGE = 32'h00000010;  // 链路状态变化中断
    localparam INT_DMA_COMPLETE = 32'h00000020; // DMA完成中断
    localparam INT_BUFFER_FULL = 32'h00000040;  // 缓冲区满中断

    always @ ( posedge clk ) begin
        if (rst) begin
            number <= 0;
            rx_packets <= 0;
            tx_packets <= 0;
            rx_bytes <= 0;
            tx_bytes <= 0;
            rx_errors <= 0;
            tx_errors <= 0;
            device_state <= 0;
            device_temperature <= 4;
            signal_strength <= 0;
            link_status <= 0;
            int_status <= 0;
            int_cause <= 0;
            int_ack <= 0;
            msix_pba <= 0;
            
            // 初始化MSI-X表
            for (int i = 0; i < 16; i++) begin
                msix_table[i] <= {32'h00000000,    // 消息地址高32位
                                  32'h00000000,    // 消息地址低32位
                                  32'h00000000,    // 消息数据
                                  32'h00000001};   // 向量控制 (已启用)
            end
        end else begin
            number          <= number + 1;
            drd_req_ctx     <= rd_req_ctx;
            drd_req_valid   <= rd_req_valid;
            dwr_valid       <= wr_valid;
            drd_req_addr    <= rd_req_addr;
            rd_rsp_ctx      <= drd_req_ctx;
            rd_rsp_valid    <= drd_req_valid;
            dwr_addr        <= wr_addr;
            dwr_data        <= wr_data;
            
            // 统计信息更新
            if (number % 997 == 0) begin
                rx_packets <= rx_packets + 1;
                rx_bytes <= rx_bytes + ((number % 1500) + 64);
                int_cause <= int_cause | INT_RX_COMPLETE;  // 触发接收完成中断
            end
            
            if (number % 1009 == 0) begin
                tx_packets <= tx_packets + 1;
                tx_bytes <= tx_bytes + ((number % 1500) + 64);
                int_cause <= int_cause | INT_TX_COMPLETE;  // 触发发送完成中断
            end
            
            if (number % 50021 == 0) begin
                rx_errors <= rx_errors + 1;
                int_cause <= int_cause | INT_RX_ERROR;  // 触发接收错误中断
            end
            
            if (number % 60037 == 0) begin
                tx_errors <= tx_errors + 1;
                int_cause <= int_cause | INT_TX_ERROR;  // 触发发送错误中断
            end
            
            // DMA中断模拟 - 周期性触发DMA完成中断
            if (number % 99 == 0) begin
                int_cause <= int_cause | INT_DMA_COMPLETE;
            end
            
            // 更新中断状态寄存器 - 根据中断原因和掩码
            int_status <= int_cause & int_mask;
            
            // 更新MSI-X PBA - 当有中断发生且对应的MSI-X表项未被屏蔽时
            if (int_cause != 0) begin
                // 设置MSI-X PBA位
                if (int_cause & INT_RX_COMPLETE) msix_pba[0] <= ~msix_table[0][0];  // 如果向量未屏蔽
                if (int_cause & INT_TX_COMPLETE) msix_pba[1] <= ~msix_table[1][0];
                if (int_cause & INT_RX_ERROR) msix_pba[2] <= ~msix_table[2][0];
                if (int_cause & INT_TX_ERROR) msix_pba[3] <= ~msix_table[3][0];
                if (int_cause & INT_LINK_CHANGE) msix_pba[4] <= ~msix_table[4][0];
                if (int_cause & INT_DMA_COMPLETE) msix_pba[5] <= ~msix_table[5][0];
                if (int_cause & INT_BUFFER_FULL) msix_pba[6] <= ~msix_table[6][0];
            end
            
            // 处理中断确认 - 如果写入了中断确认寄存器，清除相应的中断原因位
            if (dwr_valid && ({dwr_addr[31:24], dwr_addr[23:16], dwr_addr[15:08], dwr_addr[07:00]} - base_address_register) == 16'h4034) begin
                int_cause <= int_cause & ~dwr_data;  // 清除已确认的中断
                
                // 同时清除对应的MSI-X PBA位
                if (dwr_data & INT_RX_COMPLETE) msix_pba[0] <= 0;
                if (dwr_data & INT_TX_COMPLETE) msix_pba[1] <= 0;
                if (dwr_data & INT_RX_ERROR) msix_pba[2] <= 0;
                if (dwr_data & INT_TX_ERROR) msix_pba[3] <= 0;
                if (dwr_data & INT_LINK_CHANGE) msix_pba[4] <= 0;
                if (dwr_data & INT_DMA_COMPLETE) msix_pba[5] <= 0;
                if (dwr_data & INT_BUFFER_FULL) msix_pba[6] <= 0;
            end
            
            // 设备状态更新
            case (device_state)
                0: if (number > 5000) device_state <= 1;
                1: if (number % 500000 == 0) device_state <= 2;
                2: if (number % 100000 == 0) device_state <= 1;
                default: if (number % 1000000 == 0) device_state <= 0;
            endcase
            
            // 温度变化
            if (number % 10000 == 0) begin
                if (device_temperature < 4) device_temperature <= 4;
                else if (device_temperature > 12) device_temperature <= 12;
                else device_temperature <= device_temperature + ((number % 3) - 1);
            end
            
            // 信号强度变化
            if (number % 15000 == 0) begin
                if (link_status == 2) signal_strength <= 8 + (number % 8);
                else signal_strength <= number % 5;
            end
            
            // 链接状态变化 - 修改为更稳定的链接状态
            if (number < 10000) begin  // 只在初始阶段变化
                case (link_status)
                    0: if (number > 2000) link_status <= 1;
                    1: if (number > 4000) link_status <= 2;
                    default: link_status <= 2;  // 保持连接状态
                endcase
            end else begin
                link_status <= 2;  // 始终保持连接状态
            end

            if (drd_req_valid)
                case ({drd_req_addr[31:24], drd_req_addr[23:16], drd_req_addr[15:08], drd_req_addr[07:00]} - base_address_register)
                    16'h2000 : begin data_32 <= 1;  rd_rsp_data <= 32'hDEADBEEF; end // EEPROM MGIC REQ
                    16'h2200 : begin data_32 <= 2;  rd_rsp_data <= 32'hDEADBEEF; end // EEPROM SIZE REQ
                    16'h2204 : begin data_32 <= 3;  rd_rsp_data <= 32'hDEADBEEF; end // EEPROM CSUM REQ
                    16'h2208 : begin data_32 <= 4;  rd_rsp_data <= 32'hDEADBEEF; end // EEPROM VERS REQ
                    16'h220C : begin data_32 <= 5;  rd_rsp_data <= 32'hDEADBEEF; end // EEPROM ANTN REQ
                    16'h2210 : begin data_32 <= 6;  rd_rsp_data <= 32'hDEADBEEF; end // EEPROM RDMN REQ
                    16'h2218 : begin data_32 <= 7;  rd_rsp_data <= 32'hDEADBEEF; end // EEPROM MAC0 REQ
                    16'h221C : begin data_32 <= 8;  rd_rsp_data <= 32'hDEADBEEF; end // EEPROM MAC1 REQ
                    16'h2220 : begin data_32 <= 9;  rd_rsp_data <= 32'hDEADBEEF; end // EEPROM MAC2 REQ
                    16'h2224 : begin data_32 <= 10; rd_rsp_data <= 32'hDEADBEEF; end // EEPROM RXTX REQ
                    16'h2228 : begin data_32 <= 11; rd_rsp_data <= 32'hDEADBEEF; end // EEPROM ENDZ REQ
                    16'h4020 : rd_rsp_data <= 32'h001800FF; // MAC VERSION
                    16'h4028 : rd_rsp_data <= int_status;   // 返回中断状态
                    16'h4030 : rd_rsp_data <= int_mask;     // 返回中断掩码
                    16'h4034 : rd_rsp_data <= int_cause;    // 返回中断原因
                    16'h4038 : rd_rsp_data <= int_status ? 32'h00000003 : 32'h00000002; // 中断状态指示
                    16'h407C :
                    case (data_32)
                        1  : rd_rsp_data <= 32'h0000A55A; // EEPROM_MAGIC
                        2  : rd_rsp_data <= 32'h00000004; // EEPROM_SIZE
                        3  : rd_rsp_data <= 32'h0000FFFB; // EEPROM_CHECKSUM
                        4  : rd_rsp_data <= 32'h0000E00E; // EEPROM_VERSION
                        5  : rd_rsp_data <= 32'h0000E00E; // EEPROM_ANTENNA (2.4ghz, 5ghz)
                        6  : rd_rsp_data <= 32'h00000000; // EEPROM_REGDOMAIN (location)
                        7  : rd_rsp_data <= 32'h0000D3C8; // EEPROM_MAC0 (C8:D3)
                        8  :
                            begin
                                rd_rsp_data[7:0]   <= 8'hA3;
                                rd_rsp_data[15:8]  <= ((0 + (number) % (15 + 1 - 0)) << 4) | (0 + (number + 3) % (15 + 1 - 0));
                                rd_rsp_data[31:16] <= 16'h0000;
                            end
                        9  :
                            begin
                                rd_rsp_data[7:0]   <= ((0 + (number + 6) % (15 + 1 - 0)) << 4) | (0 + (number + 9) % (15 + 1 - 0));
                                rd_rsp_data[15:8]  <= ((0 + (number + 12) % (15 + 1 - 0)) << 4) | (0 + (number + 15) % (15 + 1 - 0));
                                rd_rsp_data[31:16] <= 16'h0000;
                            end
                        10 : rd_rsp_data <= 32'h00000100; // EEPROM_RXTX (00,01)
                        11 : begin rd_rsp_data <= 32'h00000000; data_32 <= 0; end
                        default : rd_rsp_data <= 32'h00000000;
                    endcase
                    16'h7000 : rd_rsp_data <= 32'h00000000; // AR_RTC_RC
                    16'h7044 : rd_rsp_data <= 32'h00000002; // AR_RTC_STATUS
                    16'h8000 : rd_rsp_data <= data_32;      // AR_STA_ID0
                    16'h806C : rd_rsp_data <= 32'h00000000; // AR_OBS_BUS_1
                    16'h9820 : rd_rsp_data <= data_32;      // AR_STA_ID0
                    16'h9860 : 
                        begin
                            // 模拟真实网卡的等待状态变化
                            if (number % 13 < 3)
                                rd_rsp_data <= 32'h00000001;
                            else if (number % 13 < 6)
                                rd_rsp_data <= 32'h00000002;
                            else
                                rd_rsp_data <= 32'h00000000;
                        end
                    16'h9C00 : 
                        begin
                            // 模拟RF状态变化
                            if (number % 17 < 5)
                                rd_rsp_data <= 32'h00000001;
                            else if (number % 17 < 10)
                                rd_rsp_data <= 32'h00000002;
                            else
                                rd_rsp_data <= 32'h00000000;
                        end
                    
                    // 统计信息寄存器 - 使用未占用的地址范围
                    16'hA000 : rd_rsp_data <= rx_packets;   // 接收数据包计数
                    16'hA004 : rd_rsp_data <= tx_packets;   // 发送数据包计数
                    16'hA008 : rd_rsp_data <= rx_bytes;     // 接收字节计数
                    16'hA00C : rd_rsp_data <= tx_bytes;     // 发送字节计数
                    16'hA010 : rd_rsp_data <= rx_errors;    // 接收错误计数
                    16'hA014 : rd_rsp_data <= tx_errors;    // 发送错误计数
                    16'hA018 : rd_rsp_data <= number[31:0]; // 运行时间计数器
                    
                    // 设备状态寄存器 - 使用未占用的地址范围
                    16'hA100 : rd_rsp_data <= {24'h0, device_state, device_temperature};  // 设备状态和温度
                    16'hA104 : rd_rsp_data <= {24'h0, signal_strength, 2'b00, link_status};  // 信号强度和链接状态
                    16'hA108 : rd_rsp_data <= 32'h00000001;  // 链接活动标志 - 始终为活动状态
                    16'hA10C : rd_rsp_data <= {8'h0, 8'h01, 8'h03, 8'h01};  // 高速能力标志
                    
                    // 添加高速链路能力寄存器
                    16'hA110 : rd_rsp_data <= 32'h00000064;  // 100Mbps能力
                    16'hA114 : rd_rsp_data <= 32'h000003E8;  // 1000Mbps能力
                    16'hA118 : rd_rsp_data <= 32'h00000001;  // 高速模式启用
                    16'hA11C : rd_rsp_data <= 32'h00000002;  // 全双工模式
                    
                    // 添加媒体类型和链路状态寄存器
                    16'hA120 : rd_rsp_data <= 32'h00000001;  // 铜缆介质
                    16'hA124 : rd_rsp_data <= 32'h00000001;  // 链路已建立
                    16'hA128 : rd_rsp_data <= 32'h00000000;  // 无错误
                    16'hA12C : rd_rsp_data <= 32'h000003E8;  // 当前速度 1000Mbps
                    
                    // 固件版本信息寄存器 - 使用未占用的地址范围
                    16'hA200 : rd_rsp_data <= 32'h02010003;  // 固件版本号: 2.1.0.3
                    16'hA204 : rd_rsp_data <= 32'h20230615;  // 固件日期: 2023/06/15
                    16'hA208 : rd_rsp_data <= 32'h41523932;  // 芯片ID "AR92" (ASCII)
                    16'hA20C : rd_rsp_data <= 32'h38370000;  // 芯片ID "87" (ASCII)
                    16'hA210 : rd_rsp_data <= 32'h44574135;  // 产品ID "DWA5" (ASCII)
                    16'hA214 : rd_rsp_data <= 32'h35360000;  // 产品ID "56" (ASCII)
                    16'hA218 : rd_rsp_data <= 32'h00000002;  // 硬件版本
                    16'hA21C : rd_rsp_data <= 32'h00000001;  // 硬件修订版本
                    
                    // MSI-X表区域 (0x0000-0x07FF)
                    // 每个表项16字节(128位)，共16个表项
                    16'h0000, 16'h0004, 16'h0008, 16'h000C: rd_rsp_data <= msix_table[0][({drd_req_addr[3:2], 5'b00000})+:32];
                    16'h0010, 16'h0014, 16'h0018, 16'h001C: rd_rsp_data <= msix_table[1][({drd_req_addr[3:2], 5'b00000})+:32];
                    16'h0020, 16'h0024, 16'h0028, 16'h002C: rd_rsp_data <= msix_table[2][({drd_req_addr[3:2], 5'b00000})+:32];
                    16'h0030, 16'h0034, 16'h0038, 16'h003C: rd_rsp_data <= msix_table[3][({drd_req_addr[3:2], 5'b00000})+:32];
                    16'h0040, 16'h0044, 16'h0048, 16'h004C: rd_rsp_data <= msix_table[4][({drd_req_addr[3:2], 5'b00000})+:32];
                    16'h0050, 16'h0054, 16'h0058, 16'h005C: rd_rsp_data <= msix_table[5][({drd_req_addr[3:2], 5'b00000})+:32];
                    16'h0060, 16'h0064, 16'h0068, 16'h006C: rd_rsp_data <= msix_table[6][({drd_req_addr[3:2], 5'b00000})+:32];
                    16'h0070, 16'h0074, 16'h0078, 16'h007C: rd_rsp_data <= msix_table[7][({drd_req_addr[3:2], 5'b00000})+:32];
                    16'h0080, 16'h0084, 16'h0088, 16'h008C: rd_rsp_data <= msix_table[8][({drd_req_addr[3:2], 5'b00000})+:32];
                    16'h0090, 16'h0094, 16'h0098, 16'h009C: rd_rsp_data <= msix_table[9][({drd_req_addr[3:2], 5'b00000})+:32];
                    16'h00A0, 16'h00A4, 16'h00A8, 16'h00AC: rd_rsp_data <= msix_table[10][({drd_req_addr[3:2], 5'b00000})+:32];
                    16'h00B0, 16'h00B4, 16'h00B8, 16'h00BC: rd_rsp_data <= msix_table[11][({drd_req_addr[3:2], 5'b00000})+:32];
                    16'h00C0, 16'h00C4, 16'h00C8, 16'h00CC: rd_rsp_data <= msix_table[12][({drd_req_addr[3:2], 5'b00000})+:32];
                    16'h00D0, 16'h00D4, 16'h00D8, 16'h00DC: rd_rsp_data <= msix_table[13][({drd_req_addr[3:2], 5'b00000})+:32];
                    16'h00E0, 16'h00E4, 16'h00E8, 16'h00EC: rd_rsp_data <= msix_table[14][({drd_req_addr[3:2], 5'b00000})+:32];
                    16'h00F0, 16'h00F4, 16'h00F8, 16'h00FC: rd_rsp_data <= msix_table[15][({drd_req_addr[3:2], 5'b00000})+:32];
                    
                    // MSI-X PBA区域 (0x0800-0x080F)
                    16'h0800: rd_rsp_data <= msix_pba;
                    16'h0804, 16'h0808, 16'h080C: rd_rsp_data <= 32'h00000000;
                    
                    default : rd_rsp_data <= 32'hDEADBEEF;  // default value: 0xDEADBEEF
                endcase
            else if (dwr_valid)
                case ({dwr_addr[31:24], dwr_addr[23:16], dwr_addr[15:08], dwr_addr[07:00]} - base_address_register)
                    16'h8000 : data_32 <= dwr_data;
                    16'h9820 : data_32 <= dwr_data;
                    16'h4030 : int_mask <= dwr_data;     // 写入中断掩码
                    16'h4034 : int_ack <= dwr_data;      // 写入中断确认
                    
                    // MSI-X表区域写入
                    16'h0000, 16'h0004, 16'h0008, 16'h000C: msix_table[0][({dwr_addr[3:2], 5'b00000})+:32] <= dwr_data;
                    16'h0010, 16'h0014, 16'h0018, 16'h001C: msix_table[1][({dwr_addr[3:2], 5'b00000})+:32] <= dwr_data;
                    16'h0020, 16'h0024, 16'h0028, 16'h002C: msix_table[2][({dwr_addr[3:2], 5'b00000})+:32] <= dwr_data;
                    16'h0030, 16'h0034, 16'h0038, 16'h003C: msix_table[3][({dwr_addr[3:2], 5'b00000})+:32] <= dwr_data;
                    16'h0040, 16'h0044, 16'h0048, 16'h004C: msix_table[4][({dwr_addr[3:2], 5'b00000})+:32] <= dwr_data;
                    16'h0050, 16'h0054, 16'h0058, 16'h005C: msix_table[5][({dwr_addr[3:2], 5'b00000})+:32] <= dwr_data;
                    16'h0060, 16'h0064, 16'h0068, 16'h006C: msix_table[6][({dwr_addr[3:2], 5'b00000})+:32] <= dwr_data;
                    16'h0070, 16'h0074, 16'h0078, 16'h007C: msix_table[7][({dwr_addr[3:2], 5'b00000})+:32] <= dwr_data;
                    16'h0080, 16'h0084, 16'h0088, 16'h008C: msix_table[8][({dwr_addr[3:2], 5'b00000})+:32] <= dwr_data;
                    16'h0090, 16'h0094, 16'h0098, 16'h009C: msix_table[9][({dwr_addr[3:2], 5'b00000})+:32] <= dwr_data;
                    16'h00A0, 16'h00A4, 16'h00A8, 16'h00AC: msix_table[10][({dwr_addr[3:2], 5'b00000})+:32] <= dwr_data;
                    16'h00B0, 16'h00B4, 16'h00B8, 16'h00BC: msix_table[11][({dwr_addr[3:2], 5'b00000})+:32] <= dwr_data;
                    16'h00C0, 16'h00C4, 16'h00C8, 16'h00CC: msix_table[12][({dwr_addr[3:2], 5'b00000})+:32] <= dwr_data;
                    16'h00D0, 16'h00D4, 16'h00D8, 16'h00DC: msix_table[13][({dwr_addr[3:2], 5'b00000})+:32] <= dwr_data;
                    16'h00E0, 16'h00E4, 16'h00E8, 16'h00EC: msix_table[14][({dwr_addr[3:2], 5'b00000})+:32] <= dwr_data;
                    16'h00F0, 16'h00F4, 16'h00F8, 16'h00FC: msix_table[15][({dwr_addr[3:2], 5'b00000})+:32] <= dwr_data;
                endcase
            else
                rd_rsp_data <= 32'hDEADBEEF;
        end
    end

endmodule

